module k_16_invsqr(input [15:0]in, input clk, output [15:0]out);
wire [4:0] ea,exponent;
reg [9:0] Rt;
assign ea=(in[14:10]-5'd15)<<1'b1;
assign exponent=5'd15-ea;
assign out={1'b0,exponent,Rt};

always @(posedge clk)
begin
if(in[9:0]<10'b0000110111) //1.053725
Rt=10'b1111001011; //0.949009587
else if(in[9:0]<10'b0001110010) //1.111895
Rt=10'b1101101001; //0.853506695
else if(in[9:0]<10'b0010110001) //1.17344
Rt=10'b1100010000; //0.766431653
else if(in[9:0]<10'b0011110010) //1.237195
Rt=10'b1011000001; //0.688809539
else if(in[9:0]<10'b0100110101) //1.302105
Rt=10'b1001111011; //0.62074628
else if(in[9:0]<10'b0101111000) //1.367345
Rt=10'b1000111111; //0.561660987
else if(in[9:0]<10'b0110111010) //1.43239
Rt=10'b1000001010; //0.510574429
else if(in[9:0]<10'b0111111100) //1.496985
Rt=10'b0111011101; //0.466358383
else if(in[9:0]<10'b1000111110) //1.561005
Rt=10'b0110110110; //0.427934043
else if(in[9:0]<10'b1001111111) //1.624395
Rt=10'b0110010011; //0.394368935
else if(in[9:0]<10'b1010111111) //1.687125
Rt=10'b0101110101; //0.36488817
else if(in[9:0]<10'b1011111111) //1.74921
Rt=10'b0101011010; //0.338851587
else if(in[9:0]<10'b1100111110) //1.81082
Rt=10'b0101000011;  //0.315705062
else if(in[9:0]<10'b1101111101) //1.87244
Rt=10'b0100101110; //0.294927743
else if(in[9:0]<10'b1110111101) //1.935005
Rt=10'b0100011010; //0.275999857
else
Rt=10'b0100001000; //0.258396608
end

endmodule