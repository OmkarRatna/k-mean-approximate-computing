module k_16_divider(input [15:0]in1,in2,input clk,en, output [15:0]out,output reg done);
reg [9:0] Rt;
reg [21:0] mul_o;
wire [5:0] exponent;
assign exponent=(in1[14:10]-in2[14:10])+4'd15;
assign out={1'b0,exponent,mul_o[20:11]};

always@(*)
begin
if(in2<10'b0000111011)				//1.05842
Rt<=10'b1111100011;	//0.971877646
else if(in2<10'b0001111011)			//1.12012
Rt<=10'b1110101100;	//0.918289501
else if(in2<10'b0010111100)			//1.184015
Rt<=10'b1101111001;	//0.868225408
else if(in2<10'b0011111111)			//1.24906
Rt<=10'b1101001001;	//0.822199295
else if(in2<10'b0101000001)			//1.314425
Rt<=10'b1100011111;	//0.780355537
else if(in2<10'b0110000100)			//1.37956
Rt<=10'b1011111000;	//0.742537964
else if(in2<10'b0111000110)			//1.444195
Rt<=10'b1011010101;	//0.708399227
else if(in2<10'b1000001000)			//1.50823
Rt<=10'b1010110101;	//0.677514351
else if(in2<10'b1001001001)			//1.571625
Rt<=10'b1010011001;	//0.649471902
else if(in2<10'b1010001001)			//1.63435
Rt<=10'b1001111110;	//0.623913827	
else if(in2<10'b1011001001)			//1.696345
Rt<=10'b1001100110;	//0.600543734
else if(in2<10'b1100000111)			//1.75755
Rt<=10'b1001010001;	//0.579116183
else if(in2<10'b1101000101)			//1.818045
Rt<=10'b1000111100;	//0.559400063
else if(in2<10'b1110000011)			//1.87812
Rt<=10'b1000101010;	//0.541148308
else if(in2<10'b1111000000)			//1.93843
Rt<=10'b1000011000:  //0.524076424
else
Rt<=10'b1000001000;	//0.507857297
end

always@(posedge clk)
begin
if(en)
	begin
		mul_o={1'b1,in1[9:0]}*{1'b0,Rt};
		done=1'b1;
	end
else
	begin
		mul_o=22'd0;
		done=1'b0;
	end
end
endmodule